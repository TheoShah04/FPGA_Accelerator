`include "vector_pkg.svh"
`include "common_defs.svh"

module sdfSphere(
    input logic clk,
    input logic rst,
    input logic valid_in,
    input vec3 p,
    input fp radius,
    output fp outputDistance,
    output logic valid_out_sphere
);
    fp vectorLength; 
    logic module_finished;

    logic q_valid_in;
    vec3  q_p;

    always_ff @ (posedge clk) begin
        q_valid_in <= valid_in;
        q_p <= p;
    end

    vec3Length calcLength(
        .clk(clk),
        .rst(rst),
        .vec(q_p),
        .valid_in(q_valid_in),
        .length(vectorLength),
        .valid_out(module_finished)
    );
    assign outputDistance = vectorLength - radius;
    assign valid_out_sphere = module_finished;

endmodule
